module text_4_bit;
reg[3:0] A;
reg[3:0] B;
reg C0;
wire [3:0] S;
wire C4;
four_bit_adder dut(A,B,C0,S,C4);
initial
begin
        A=4'B0011; B=4'B0011; C0=1'B0;
#10; A=4'B0000; B=4'B0000; C0=1'B1;
#10; A=4'B0001; B=4'B0001; C0=1'B0;
#10; A=4'B0001; B=4'B0001; C0=1'B1;
#10; A=4'B0010; B=4'B0010; C0=1'B0;
#10; A=4'B0010; B=4'B0010; C0=1'B1;
#10; A=4'B0011; B=4'B0011; C0=1'B0;
#10; A=4'B0011; B=4'B0011; C0=1'B1;
#10; A=4'B0100; B=4'B0100; C0=1'B0;
#10; A=4'B0100; B=4'B0100; C0=1'B1;
#10; A=4'B0101; B=4'B0101; C0=1'B0;
#10; A=4'B0101; B=4'B0101; C0=1'B1;
#10; A=4'B0110; B=4'B0110; C0=1'B0;
#10; A=4'B0110; B=4'B0110; C0=1'B1;
#10; A=4'B0111; B=4'B0111; C0=1'B0;
#10; A=4'B0111; B=4'B0111; C0=1'B1;
#10; A=4'B1000; B=4'B1000; C0=1'B0;
#10; A=4'B1000; B=4'B1000; C0=1'B1;
#10; A=4'B1001; B=4'B1001; C0=1'B0;
#10; A=4'B1001; B=4'B1001; C0=1'B1;
#10; A=4'B1010; B=4'B1010; C0=1'B0;
#10; A=4'B1010; B=4'B1010; C0=1'B1;
#10; A=4'B1011; B=4'B1011; C0=1'B0;
#10; A=4'B1011; B=4'B1011; C0=1'B1;
#10; A=4'B1100; B=4'B1100; C0=1'B0;
#10; A=4'B1100; B=4'B1100; C0=1'B1;
#10; A=4'B1101; B=4'B1101; C0=1'B0;
#10; A=4'B1101; B=4'B1101; C0=1'B1;
#10; A=4'B1110; B=4'B1110; C0=1'B0;
#10; A=4'B1110; B=4'B1110; C0=1'B1;
#10; A=4'B1111; B=4'B1111; C0=1'B0;
#10; A=4'B1111; B=4'B1111; C0=1'B1;
#10; A=4'B0001; B=4'B0001; C0=1'B0;

end
initial
#50 $finish;
endmodule



